module control(opcode, RegDst, Branch, ALUSrc, MemWrite, MemRead, MentoReg);
	input wire [5:0] opcode;
	output wire RegDst;
	output wire Branch;
	output wire ALUSrc;
	output wire MemWrite;
	output wire MemRead;
	output wire MentoReg;

	
	//seria a descricao do circuito
	
endmodule 