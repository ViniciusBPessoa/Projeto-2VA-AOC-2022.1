module control(opcode, RegDst, Branch, ALUSrc, MemWrite, MemRead, MentoReg, ALUOp, MenWrite);
	input wire [5:0] opcode;
	output wire RegDst;
	output wire Branch;
	output wire ALUSrc;
	output wire MemWrite;
	output wire MemRead;
	output wire MentoReg;
	output wire MenWrite;
	output wire [3:0] ALUOp;

	
	//seria a descricao do circuito
	
endmodule 